module ALU();

endmodule
