module Decoder
